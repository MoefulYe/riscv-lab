module InstMem(
    input clk,
    input [31:0] addr, //addr[7:2]
    output [31:0] inst
);

endmodule