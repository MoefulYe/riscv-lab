`include "../03-ALU/ALU.v"
`include "../04-reg-heap/RegHeap.v"
`include "../07-inst-fetch-decode/ProgramCounter.v"
`include "../07-inst-fetch-decode/InstDecoder1.v"

module CU (

);
endmodule

module CPUimplRIU(
    input clk,
    input rst,

);
endmodule